LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY TestBCDCount2_G02 IS
	PORT (KEY					: IN STD_LOGIC_VECTOR (1 DOWNTO 0);
			SW						: IN STD_LOGIC_VECTOR(0 DOWNTO 0);
			LEDR					: OUT STD_LOGIC_VECTOR(7 DOWNTO 0));
END TestBCDCount2_G02;

ARCHITECTURE Behaviour OF TestBCDCount2_G02 IS
COMPONENT BCDCount2_G02 IS
	PORT (clear, enable, clock		: IN STD_LOGIC;
			BCD0, BCD1					: OUT STD_LOGIC_VECTOR(3 DOWNTO 0));
END COMPONENT;
BEGIN
U1: BCDCount2_G02 PORT MAP (NOT(KEY(0)), SW(0), NOT(KEY(1)), LEDR(3 DOWNTO 0), LEDR(7 DOWNTO 4));
END Behaviour;
